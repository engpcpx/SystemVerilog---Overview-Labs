/*
    A testbench is provided in the scale_mux_test.sv file. Simulate the testbench
    and MUX design.
    You should see the following results:
    0ns in_a=00 in_b=00 sel_a=0 out=00
    1ns in_a=00 in_b=00 sel_a=1 out=00
    2ns in_a=00 in_b=ff sel_a=0 out=ff
    3ns in_a=00 in_b=ff sel_a=1 out=00
    4ns in_a=ff in_b=00 sel_a=0 out=00
    5ns in_a=ff in_b=00 sel_a=1 out=ff
    6ns in_a=ff in_b=ff sel_a=0 out=ff
    7ns in_a=ff in_b=ff sel_a=1 out=ff
    MUX TEST PASSED
*/

module scale_mux_test();


endmodule