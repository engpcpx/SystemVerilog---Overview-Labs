/*
    Lab 1 - Modeling a Simple Register Testbech


*/
'timescale 1ns/1ps
module register_tb();

