


module register (
    
);